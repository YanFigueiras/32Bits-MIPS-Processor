LIBRARY IEEE;
use ieee.std_logic_1164.all;

Entity leftShift2 is
port (
entrada: in std_logic_vector (31 downto 0);
saida: out std_logic_vector (31 downto 0)
);
end leftShift2;

architecture Leftshift2 of leftShift2 is
begin
saida <= entrada(29 downto 0) & "00"; 
end Leftshift2;